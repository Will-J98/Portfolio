<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-7.81444,1.42076,149.011,-77.5542</PageViewport>
<gate>
<ID>2</ID>
<type>DD_KEYPAD_HEX</type>
<position>11.5,-11.5</position>
<output>
<ID>OUT_0</ID>11 </output>
<output>
<ID>OUT_1</ID>10 </output>
<output>
<ID>OUT_2</ID>8 </output>
<output>
<ID>OUT_3</ID>9 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 14</lparam></gate>
<gate>
<ID>4</ID>
<type>DD_KEYPAD_HEX</type>
<position>1.5,-65</position>
<output>
<ID>OUT_0</ID>83 </output>
<output>
<ID>OUT_1</ID>82 </output>
<output>
<ID>OUT_2</ID>81 </output>
<output>
<ID>OUT_3</ID>80 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 9</lparam></gate>
<gate>
<ID>6</ID>
<type>BA_DECODER_2x4</type>
<position>23,-9.5</position>
<input>
<ID>ENABLE</ID>7 </input>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT_0</ID>20 </output>
<output>
<ID>OUT_1</ID>36 </output>
<output>
<ID>OUT_2</ID>22 </output>
<output>
<ID>OUT_3</ID>23 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8</ID>
<type>BA_DECODER_2x4</type>
<position>23.5,-18</position>
<input>
<ID>ENABLE</ID>12 </input>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT_1</ID>47 </output>
<output>
<ID>OUT_2</ID>46 </output>
<output>
<ID>OUT_3</ID>45 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>12</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>25,-58</position>
<input>
<ID>ENABLE_0</ID>20 </input>
<input>
<ID>IN_0</ID>87 </input>
<input>
<ID>IN_1</ID>88 </input>
<input>
<ID>IN_2</ID>85 </input>
<input>
<ID>IN_3</ID>84 </input>
<output>
<ID>OUT_0</ID>31 </output>
<output>
<ID>OUT_1</ID>30 </output>
<output>
<ID>OUT_2</ID>29 </output>
<output>
<ID>OUT_3</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_REGISTER4</type>
<position>34,-38</position>
<input>
<ID>IN_0</ID>56 </input>
<input>
<ID>IN_1</ID>55 </input>
<input>
<ID>IN_2</ID>54 </input>
<input>
<ID>IN_3</ID>52 </input>
<output>
<ID>OUT_0</ID>40 </output>
<output>
<ID>OUT_1</ID>39 </output>
<output>
<ID>OUT_2</ID>38 </output>
<output>
<ID>OUT_3</ID>37 </output>
<input>
<ID>clear</ID>13 </input>
<input>
<ID>clock</ID>25 </input>
<input>
<ID>count_enable</ID>1 </input>
<input>
<ID>count_up</ID>2 </input>
<input>
<ID>load</ID>45 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_REGISTER4</type>
<position>66.5,-41</position>
<input>
<ID>IN_0</ID>70 </input>
<input>
<ID>IN_1</ID>69 </input>
<input>
<ID>IN_2</ID>67 </input>
<input>
<ID>IN_3</ID>66 </input>
<output>
<ID>OUT_0</ID>35 </output>
<output>
<ID>OUT_1</ID>34 </output>
<output>
<ID>OUT_2</ID>33 </output>
<output>
<ID>OUT_3</ID>32 </output>
<input>
<ID>clear</ID>14 </input>
<input>
<ID>clock</ID>27 </input>
<input>
<ID>count_enable</ID>3 </input>
<input>
<ID>count_up</ID>4 </input>
<input>
<ID>load</ID>46 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_REGISTER4</type>
<position>84,-23.5</position>
<input>
<ID>IN_0</ID>65 </input>
<input>
<ID>IN_1</ID>64 </input>
<input>
<ID>IN_2</ID>62 </input>
<input>
<ID>IN_3</ID>61 </input>
<output>
<ID>OUT_0</ID>51 </output>
<output>
<ID>OUT_1</ID>50 </output>
<output>
<ID>OUT_2</ID>49 </output>
<output>
<ID>OUT_3</ID>48 </output>
<input>
<ID>clear</ID>15 </input>
<input>
<ID>clock</ID>26 </input>
<input>
<ID>count_enable</ID>6 </input>
<input>
<ID>count_up</ID>5 </input>
<input>
<ID>load</ID>47 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>20</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>103,-57</position>
<input>
<ID>IN_0</ID>44 </input>
<input>
<ID>IN_1</ID>43 </input>
<input>
<ID>IN_2</ID>42 </input>
<input>
<ID>IN_3</ID>41 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>22</ID>
<type>FF_GND</type>
<position>34.5,-30.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>24</ID>
<type>FF_GND</type>
<position>33.5,-30.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>26</ID>
<type>EE_VDD</type>
<position>17,-8</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>27</ID>
<type>FF_GND</type>
<position>65.5,-32</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>28</ID>
<type>FF_GND</type>
<position>85,-14.5</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>29</ID>
<type>FF_GND</type>
<position>66.5,-34</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>30</ID>
<type>FF_GND</type>
<position>84,-16</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>32</ID>
<type>EE_VDD</type>
<position>20,-14.5</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>34</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>43,-37.5</position>
<input>
<ID>ENABLE_0</ID>36 </input>
<input>
<ID>IN_0</ID>40 </input>
<input>
<ID>IN_1</ID>39 </input>
<input>
<ID>IN_2</ID>38 </input>
<input>
<ID>IN_3</ID>37 </input>
<output>
<ID>OUT_0</ID>60 </output>
<output>
<ID>OUT_1</ID>59 </output>
<output>
<ID>OUT_2</ID>58 </output>
<output>
<ID>OUT_3</ID>57 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>36</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>74,-40.5</position>
<input>
<ID>ENABLE_0</ID>22 </input>
<input>
<ID>IN_0</ID>35 </input>
<input>
<ID>IN_1</ID>34 </input>
<input>
<ID>IN_2</ID>33 </input>
<input>
<ID>IN_3</ID>32 </input>
<output>
<ID>OUT_0</ID>76 </output>
<output>
<ID>OUT_1</ID>77 </output>
<output>
<ID>OUT_2</ID>78 </output>
<output>
<ID>OUT_3</ID>79 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>38</ID>
<type>FF_GND</type>
<position>34.5,-45</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>40</ID>
<type>FF_GND</type>
<position>66.5,-47.5</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>42</ID>
<type>FF_GND</type>
<position>85,-29.5</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>44</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>92,-23</position>
<input>
<ID>ENABLE_0</ID>23 </input>
<input>
<ID>IN_0</ID>51 </input>
<input>
<ID>IN_1</ID>50 </input>
<input>
<ID>IN_2</ID>49 </input>
<input>
<ID>IN_3</ID>48 </input>
<output>
<ID>OUT_0</ID>72 </output>
<output>
<ID>OUT_1</ID>73 </output>
<output>
<ID>OUT_2</ID>74 </output>
<output>
<ID>OUT_3</ID>75 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>46</ID>
<type>AA_TOGGLE</type>
<position>16,-72</position>
<output>
<ID>OUT_0</ID>24 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>48</ID>
<type>DE_TO</type>
<position>27.5,-69</position>
<input>
<ID>IN_0</ID>24 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Clock</lparam></gate>
<gate>
<ID>50</ID>
<type>DA_FROM</type>
<position>32.5,-47</position>
<input>
<ID>IN_0</ID>25 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Clock</lparam></gate>
<gate>
<ID>51</ID>
<type>DA_FROM</type>
<position>64.5,-48</position>
<input>
<ID>IN_0</ID>27 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Clock</lparam></gate>
<gate>
<ID>52</ID>
<type>DA_FROM</type>
<position>83,-30.5</position>
<input>
<ID>IN_0</ID>26 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Clock</lparam></gate>
<gate>
<ID>54</ID>
<type>DE_TO</type>
<position>34.5,-55.5</position>
<input>
<ID>IN_0</ID>28 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>56</ID>
<type>DE_TO</type>
<position>41,-57.5</position>
<input>
<ID>IN_0</ID>29 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>58</ID>
<type>DE_TO</type>
<position>47,-60</position>
<input>
<ID>IN_0</ID>30 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>60</ID>
<type>DE_TO</type>
<position>50.5,-63</position>
<input>
<ID>IN_0</ID>31 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>62</ID>
<type>DA_FROM</type>
<position>79,-53</position>
<input>
<ID>IN_0</ID>41 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>64</ID>
<type>DA_FROM</type>
<position>86,-55.5</position>
<input>
<ID>IN_0</ID>42 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>66</ID>
<type>DA_FROM</type>
<position>90,-58.5</position>
<input>
<ID>IN_0</ID>43 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>68</ID>
<type>DA_FROM</type>
<position>92.5,-62</position>
<input>
<ID>IN_0</ID>44 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>69</ID>
<type>DA_FROM</type>
<position>20.5,-36</position>
<input>
<ID>IN_0</ID>52 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>70</ID>
<type>DA_FROM</type>
<position>20.5,-38.5</position>
<input>
<ID>IN_0</ID>54 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>71</ID>
<type>DA_FROM</type>
<position>19.5,-41.5</position>
<input>
<ID>IN_0</ID>55 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>73</ID>
<type>DA_FROM</type>
<position>20,-45</position>
<input>
<ID>IN_0</ID>56 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>74</ID>
<type>DE_TO</type>
<position>49.5,-43</position>
<input>
<ID>IN_0</ID>57 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>75</ID>
<type>DE_TO</type>
<position>47,-43</position>
<input>
<ID>IN_0</ID>58 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>76</ID>
<type>DE_TO</type>
<position>44.5,-43</position>
<input>
<ID>IN_0</ID>59 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>77</ID>
<type>DE_TO</type>
<position>41.5,-43</position>
<input>
<ID>IN_0</ID>60 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>78</ID>
<type>DA_FROM</type>
<position>58,-37</position>
<input>
<ID>IN_0</ID>66 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>79</ID>
<type>DA_FROM</type>
<position>58,-39.5</position>
<input>
<ID>IN_0</ID>67 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>80</ID>
<type>DA_FROM</type>
<position>57.5,-42.5</position>
<input>
<ID>IN_0</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>81</ID>
<type>DA_FROM</type>
<position>57.5,-46</position>
<input>
<ID>IN_0</ID>70 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>82</ID>
<type>DA_FROM</type>
<position>76,-21</position>
<input>
<ID>IN_0</ID>61 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>83</ID>
<type>DA_FROM</type>
<position>76,-23.5</position>
<input>
<ID>IN_0</ID>62 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>84</ID>
<type>DA_FROM</type>
<position>75,-26.5</position>
<input>
<ID>IN_0</ID>64 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>85</ID>
<type>DA_FROM</type>
<position>75.5,-30</position>
<input>
<ID>IN_0</ID>65 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>86</ID>
<type>DE_TO</type>
<position>85.5,-44.5</position>
<input>
<ID>IN_0</ID>79 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>87</ID>
<type>DE_TO</type>
<position>83,-44.5</position>
<input>
<ID>IN_0</ID>78 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>88</ID>
<type>DE_TO</type>
<position>80.5,-44.5</position>
<input>
<ID>IN_0</ID>77 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>89</ID>
<type>DE_TO</type>
<position>77.5,-44.5</position>
<input>
<ID>IN_0</ID>76 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>90</ID>
<type>DE_TO</type>
<position>104.5,-27.5</position>
<input>
<ID>IN_0</ID>75 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>91</ID>
<type>DE_TO</type>
<position>102,-27.5</position>
<input>
<ID>IN_0</ID>74 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>92</ID>
<type>DE_TO</type>
<position>99.5,-27.5</position>
<input>
<ID>IN_0</ID>73 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>93</ID>
<type>DE_TO</type>
<position>96.5,-27.5</position>
<input>
<ID>IN_0</ID>72 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>95</ID>
<type>AA_RAM_4x4</type>
<position>16.5,-57.5</position>
<input>
<ID>ADDRESS_0</ID>83 </input>
<input>
<ID>ADDRESS_1</ID>82 </input>
<input>
<ID>ADDRESS_2</ID>81 </input>
<input>
<ID>ADDRESS_3</ID>80 </input>
<input>
<ID>DATA_IN_0</ID>84 </input>
<input>
<ID>DATA_IN_1</ID>85 </input>
<input>
<ID>DATA_IN_2</ID>88 </input>
<input>
<ID>DATA_IN_3</ID>87 </input>
<output>
<ID>DATA_OUT_0</ID>84 </output>
<output>
<ID>DATA_OUT_1</ID>85 </output>
<output>
<ID>DATA_OUT_2</ID>88 </output>
<output>
<ID>DATA_OUT_3</ID>87 </output>
<gparam>angle 90</gparam>
<lparam>ADDRESS_BITS 4</lparam>
<lparam>DATA_BITS 4</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>13</ID>
<points>34,-33,34,-31.5</points>
<connection>
<GID>14</GID>
<name>count_enable</name></connection>
<intersection>-31.5 16</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>33.5,-31.5,34,-31.5</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>34 13</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-33,35,-31.5</points>
<connection>
<GID>14</GID>
<name>count_up</name></connection>
<intersection>-31.5 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>34.5,-31.5,35,-31.5</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-36,66.5,-33</points>
<connection>
<GID>16</GID>
<name>count_enable</name></connection>
<intersection>-33 12</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>65.5,-33,66.5,-33</points>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection>
<intersection>66.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>66.5,-35,67.5,-35</points>
<connection>
<GID>29</GID>
<name>OUT_0</name></connection>
<intersection>67.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>67.5,-36,67.5,-35</points>
<connection>
<GID>16</GID>
<name>count_up</name></connection>
<intersection>-35 6</intersection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,-18.5,85,-15.5</points>
<connection>
<GID>18</GID>
<name>count_up</name></connection>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,-18.5,84,-17</points>
<connection>
<GID>18</GID>
<name>count_enable</name></connection>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>18,-8,20,-8</points>
<connection>
<GID>6</GID>
<name>ENABLE</name></connection>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-10.5,20,-10.5</points>
<connection>
<GID>2</GID>
<name>OUT_2</name></connection>
<intersection>20 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>20,-11,20,-10.5</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>-10.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-8.5,20,-8.5</points>
<connection>
<GID>2</GID>
<name>OUT_3</name></connection>
<intersection>20 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>20,-10,20,-8.5</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>-8.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18.5,-18.5,18.5,-12.5</points>
<intersection>-18.5 1</intersection>
<intersection>-12.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18.5,-18.5,20.5,-18.5</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<intersection>18.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16.5,-12.5,18.5,-12.5</points>
<connection>
<GID>2</GID>
<name>OUT_1</name></connection>
<intersection>18.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,-19.5,17.5,-14.5</points>
<intersection>-19.5 1</intersection>
<intersection>-14.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,-19.5,20.5,-19.5</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16.5,-14.5,17.5,-14.5</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>17.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20,-16.5,20,-15.5</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20,-16.5,20.5,-16.5</points>
<connection>
<GID>8</GID>
<name>ENABLE</name></connection>
<intersection>20 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-44,35,-42</points>
<connection>
<GID>14</GID>
<name>clear</name></connection>
<intersection>-44 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>34.5,-44,35,-44</points>
<connection>
<GID>38</GID>
<name>OUT_0</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>66.5,-46.5,67.5,-46.5</points>
<connection>
<GID>40</GID>
<name>OUT_0</name></connection>
<intersection>67.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>67.5,-46.5,67.5,-45</points>
<connection>
<GID>16</GID>
<name>clear</name></connection>
<intersection>-46.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,-28.5,85,-27.5</points>
<connection>
<GID>42</GID>
<name>OUT_0</name></connection>
<connection>
<GID>18</GID>
<name>clear</name></connection></vsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-51.5,27.5,-11</points>
<intersection>-51.5 3</intersection>
<intersection>-11 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>26,-11,27.5,-11</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>25,-51.5,27.5,-51.5</points>
<intersection>25 4</intersection>
<intersection>27.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>25,-55,25,-51.5</points>
<connection>
<GID>12</GID>
<name>ENABLE_0</name></connection>
<intersection>-51.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74,-37.5,74,-9</points>
<connection>
<GID>36</GID>
<name>ENABLE_0</name></connection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-9,74,-9</points>
<connection>
<GID>6</GID>
<name>OUT_2</name></connection>
<intersection>74 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92,-20,92,-8</points>
<connection>
<GID>44</GID>
<name>ENABLE_0</name></connection>
<intersection>-8 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-8,92,-8</points>
<connection>
<GID>6</GID>
<name>OUT_3</name></connection>
<intersection>92 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17.5,-70.5,25.5,-70.5</points>
<intersection>17.5 15</intersection>
<intersection>25.5 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>25.5,-70.5,25.5,-69</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>-70.5 1</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>17.5,-72,17.5,-70.5</points>
<intersection>-72 16</intersection>
<intersection>-70.5 1</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>17.5,-72,18,-72</points>
<connection>
<GID>46</GID>
<name>OUT_0</name></connection>
<intersection>17.5 15</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-45,33,-42</points>
<connection>
<GID>14</GID>
<name>clock</name></connection>
<intersection>-45 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>32.5,-45,33,-45</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>33 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83,-28.5,83,-27.5</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<connection>
<GID>18</GID>
<name>clock</name></connection></vsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>64.5,-46,65.5,-46</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>65.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>65.5,-46,65.5,-45</points>
<connection>
<GID>16</GID>
<name>clock</name></connection>
<intersection>-46 3</intersection></vsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27,-55.5,32.5,-55.5</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>27 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>27,-56.5,27,-55.5</points>
<connection>
<GID>12</GID>
<name>OUT_3</name></connection>
<intersection>-55.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27,-57.5,39,-57.5</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>27 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>27,-57.5,27,-57.5</points>
<connection>
<GID>12</GID>
<name>OUT_2</name></connection>
<intersection>-57.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-60,35,-58.5</points>
<intersection>-60 1</intersection>
<intersection>-58.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-60,45,-60</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-58.5,35,-58.5</points>
<connection>
<GID>12</GID>
<name>OUT_1</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-63,34,-59.5</points>
<intersection>-63 1</intersection>
<intersection>-59.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-63,48.5,-63</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-59.5,34,-59.5</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70.5,-39,72,-39</points>
<connection>
<GID>16</GID>
<name>OUT_3</name></connection>
<connection>
<GID>36</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70.5,-40,72,-40</points>
<connection>
<GID>16</GID>
<name>OUT_2</name></connection>
<connection>
<GID>36</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70.5,-41,72,-41</points>
<connection>
<GID>16</GID>
<name>OUT_1</name></connection>
<connection>
<GID>36</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70.5,-42,72,-42</points>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<connection>
<GID>36</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43,-34.5,43,-10</points>
<connection>
<GID>34</GID>
<name>ENABLE_0</name></connection>
<intersection>-10 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-10,43,-10</points>
<connection>
<GID>6</GID>
<name>OUT_1</name></connection>
<intersection>43 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-36,41,-36</points>
<connection>
<GID>34</GID>
<name>IN_3</name></connection>
<connection>
<GID>14</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-37,41,-37</points>
<connection>
<GID>34</GID>
<name>IN_2</name></connection>
<connection>
<GID>14</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-38,41,-38</points>
<connection>
<GID>34</GID>
<name>IN_1</name></connection>
<connection>
<GID>14</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-39,41,-39</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>81,-53,100,-53</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<intersection>100 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>100,-55,100,-53</points>
<connection>
<GID>20</GID>
<name>IN_3</name></connection>
<intersection>-53 1</intersection></vsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>88,-55.5,100,-55.5</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<intersection>100 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>100,-56,100,-55.5</points>
<connection>
<GID>20</GID>
<name>IN_2</name></connection>
<intersection>-55.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92,-58.5,92,-57</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>-57 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>92,-57,100,-57</points>
<connection>
<GID>20</GID>
<name>IN_1</name></connection>
<intersection>92 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93.5,-62,93.5,-58</points>
<intersection>-62 2</intersection>
<intersection>-58 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>93.5,-58,100,-58</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>93.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>93.5,-62,94.5,-62</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<intersection>93.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-33,33,-16.5</points>
<connection>
<GID>14</GID>
<name>load</name></connection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-16.5,33,-16.5</points>
<connection>
<GID>8</GID>
<name>OUT_3</name></connection>
<intersection>33 0</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65.5,-36,65.5,-17.5</points>
<connection>
<GID>16</GID>
<name>load</name></connection>
<intersection>-17.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-17.5,65.5,-17.5</points>
<connection>
<GID>8</GID>
<name>OUT_2</name></connection>
<intersection>65.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-18.5,83,-18.5</points>
<connection>
<GID>18</GID>
<name>load</name></connection>
<connection>
<GID>8</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>88,-21.5,90,-21.5</points>
<connection>
<GID>44</GID>
<name>IN_3</name></connection>
<connection>
<GID>18</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>88,-22.5,90,-22.5</points>
<connection>
<GID>44</GID>
<name>IN_2</name></connection>
<connection>
<GID>18</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>88,-23.5,90,-23.5</points>
<connection>
<GID>44</GID>
<name>IN_1</name></connection>
<connection>
<GID>18</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>88,-24.5,90,-24.5</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22.5,-36,30,-36</points>
<connection>
<GID>14</GID>
<name>IN_3</name></connection>
<connection>
<GID>69</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-38.5,26,-37</points>
<intersection>-38.5 2</intersection>
<intersection>-37 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-37,30,-37</points>
<connection>
<GID>14</GID>
<name>IN_2</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22.5,-38.5,26,-38.5</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>26 0</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-41.5,26.5,-38</points>
<intersection>-41.5 2</intersection>
<intersection>-38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-38,30,-38</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21.5,-41.5,26.5,-41.5</points>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<intersection>26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-45,27,-39</points>
<intersection>-45 2</intersection>
<intersection>-39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,-39,30,-39</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22,-45,27,-45</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-41,49.5,-36</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>-36 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,-36,49.5,-36</points>
<connection>
<GID>34</GID>
<name>OUT_3</name></connection>
<intersection>49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-41,47,-37</points>
<connection>
<GID>75</GID>
<name>IN_0</name></connection>
<intersection>-37 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,-37,47,-37</points>
<connection>
<GID>34</GID>
<name>OUT_2</name></connection>
<intersection>47 0</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44.5,-41,44.5,-38</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<intersection>-38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44.5,-38,45,-38</points>
<connection>
<GID>34</GID>
<name>OUT_1</name></connection>
<intersection>44.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46.5,-41.5,46.5,-39</points>
<intersection>-41.5 2</intersection>
<intersection>-39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,-39,46.5,-39</points>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection>
<intersection>46.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>41.5,-41.5,46.5,-41.5</points>
<intersection>41.5 3</intersection>
<intersection>46.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>41.5,-41.5,41.5,-41</points>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<intersection>-41.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79,-21.5,79,-21</points>
<intersection>-21.5 1</intersection>
<intersection>-21 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>79,-21.5,80,-21.5</points>
<connection>
<GID>18</GID>
<name>IN_3</name></connection>
<intersection>79 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>78,-21,79,-21</points>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<intersection>79 0</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79,-23.5,79,-22.5</points>
<intersection>-23.5 2</intersection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>79,-22.5,80,-22.5</points>
<connection>
<GID>18</GID>
<name>IN_2</name></connection>
<intersection>79 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>78,-23.5,79,-23.5</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<intersection>79 0</intersection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78.5,-26.5,78.5,-23.5</points>
<intersection>-26.5 2</intersection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>78.5,-23.5,80,-23.5</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<intersection>78.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77,-26.5,78.5,-26.5</points>
<connection>
<GID>84</GID>
<name>IN_0</name></connection>
<intersection>78.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78.5,-30,78.5,-24.5</points>
<intersection>-30 2</intersection>
<intersection>-24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>78.5,-24.5,80,-24.5</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>78.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77.5,-30,78.5,-30</points>
<connection>
<GID>85</GID>
<name>IN_0</name></connection>
<intersection>78.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-39,60.5,-37</points>
<intersection>-39 1</intersection>
<intersection>-37 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60.5,-39,62.5,-39</points>
<connection>
<GID>16</GID>
<name>IN_3</name></connection>
<intersection>60.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>60,-37,60.5,-37</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<intersection>60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-40,60.5,-39.5</points>
<intersection>-40 1</intersection>
<intersection>-39.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60.5,-40,62.5,-40</points>
<connection>
<GID>16</GID>
<name>IN_2</name></connection>
<intersection>60.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>60,-39.5,60.5,-39.5</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61,-42.5,61,-41</points>
<intersection>-42.5 2</intersection>
<intersection>-41 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61,-41,62.5,-41</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<intersection>61 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>59.5,-42.5,61,-42.5</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<intersection>61 0</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61,-46,61,-42</points>
<intersection>-46 2</intersection>
<intersection>-42 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61,-42,62.5,-42</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>61 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>59.5,-46,61,-46</points>
<connection>
<GID>81</GID>
<name>IN_0</name></connection>
<intersection>61 0</intersection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96.5,-25.5,96.5,-24.5</points>
<connection>
<GID>93</GID>
<name>IN_0</name></connection>
<intersection>-24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>94,-24.5,96.5,-24.5</points>
<connection>
<GID>44</GID>
<name>OUT_0</name></connection>
<intersection>96.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99.5,-25.5,99.5,-23.5</points>
<connection>
<GID>92</GID>
<name>IN_0</name></connection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>94,-23.5,99.5,-23.5</points>
<connection>
<GID>44</GID>
<name>OUT_1</name></connection>
<intersection>99.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,-25.5,102,-22.5</points>
<connection>
<GID>91</GID>
<name>IN_0</name></connection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>94,-22.5,102,-22.5</points>
<connection>
<GID>44</GID>
<name>OUT_2</name></connection>
<intersection>102 0</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-25.5,104.5,-21.5</points>
<connection>
<GID>90</GID>
<name>IN_0</name></connection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>94,-21.5,104.5,-21.5</points>
<connection>
<GID>44</GID>
<name>OUT_3</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-42.5,77.5,-42</points>
<connection>
<GID>89</GID>
<name>IN_0</name></connection>
<intersection>-42 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76,-42,77.5,-42</points>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection>
<intersection>77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80.5,-42.5,80.5,-41</points>
<connection>
<GID>88</GID>
<name>IN_0</name></connection>
<intersection>-41 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76,-41,80.5,-41</points>
<connection>
<GID>36</GID>
<name>OUT_1</name></connection>
<intersection>80.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83,-42.5,83,-40</points>
<connection>
<GID>87</GID>
<name>IN_0</name></connection>
<intersection>-40 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76,-40,83,-40</points>
<connection>
<GID>36</GID>
<name>OUT_2</name></connection>
<intersection>83 0</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85.5,-42.5,85.5,-39</points>
<connection>
<GID>86</GID>
<name>IN_0</name></connection>
<intersection>-39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76,-39,85.5,-39</points>
<connection>
<GID>36</GID>
<name>OUT_3</name></connection>
<intersection>85.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>6.5,-62,15,-62</points>
<connection>
<GID>4</GID>
<name>OUT_3</name></connection>
<intersection>15 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>15,-62.5,15,-62</points>
<connection>
<GID>95</GID>
<name>ADDRESS_3</name></connection>
<intersection>-62 1</intersection></vsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,-64,16,-62.5</points>
<connection>
<GID>95</GID>
<name>ADDRESS_2</name></connection>
<intersection>-64 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>6.5,-64,16,-64</points>
<connection>
<GID>4</GID>
<name>OUT_2</name></connection>
<intersection>16 0</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,-66,17,-62.5</points>
<connection>
<GID>95</GID>
<name>ADDRESS_1</name></connection>
<intersection>-66 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>6.5,-66,17,-66</points>
<connection>
<GID>4</GID>
<name>OUT_1</name></connection>
<intersection>17 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-68,18,-62.5</points>
<connection>
<GID>95</GID>
<name>ADDRESS_0</name></connection>
<intersection>-68 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>6.5,-68,18,-68</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,-56.5,22,-56</points>
<intersection>-56.5 1</intersection>
<intersection>-56 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22,-56.5,23,-56.5</points>
<connection>
<GID>12</GID>
<name>IN_3</name></connection>
<intersection>22 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21.5,-56,22,-56</points>
<connection>
<GID>95</GID>
<name>DATA_OUT_0</name></connection>
<connection>
<GID>95</GID>
<name>DATA_IN_0</name></connection>
<intersection>22 0</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,-57.5,22,-57</points>
<intersection>-57.5 1</intersection>
<intersection>-57 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22,-57.5,23,-57.5</points>
<connection>
<GID>12</GID>
<name>IN_2</name></connection>
<intersection>22 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21.5,-57,22,-57</points>
<connection>
<GID>95</GID>
<name>DATA_OUT_1</name></connection>
<connection>
<GID>95</GID>
<name>DATA_IN_1</name></connection>
<intersection>22 0</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,-59.5,22,-59</points>
<intersection>-59.5 1</intersection>
<intersection>-59 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22,-59.5,23,-59.5</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>22 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21.5,-59,22,-59</points>
<connection>
<GID>95</GID>
<name>DATA_OUT_3</name></connection>
<connection>
<GID>95</GID>
<name>DATA_IN_3</name></connection>
<intersection>22 0</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,-58.5,22,-58</points>
<intersection>-58.5 1</intersection>
<intersection>-58 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22,-58.5,23,-58.5</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<intersection>22 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21.5,-58,22,-58</points>
<connection>
<GID>95</GID>
<name>DATA_OUT_2</name></connection>
<connection>
<GID>95</GID>
<name>DATA_IN_2</name></connection>
<intersection>22 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 1>
<page 2>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 2>
<page 3>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 3>
<page 4>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 4>
<page 5>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 5>
<page 6>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 6>
<page 7>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 7>
<page 8>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 8>
<page 9>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 9></circuit>